library ieee;
    use ieee.std_logic_1164.all;


package array_pkg is

    type slv_array_t is array (natural range <>) of std_logic_vector(31 downto 0); 
    
end package array_pkg;


package body array_pkg is

end package body array_pkg;