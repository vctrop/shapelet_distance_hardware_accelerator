library ieee;
    use ieee.std_logic_1164.all;


package AdderTreePKG is
	
	type slv_vector is array(natural range <>) of std_logic_vector(31 downto 0);

end package AdderTreePKG;


package body AdderTreePKG is

end package body AdderTreePKG;