library ieee;
    use ieee.std_logic_1164.all;


package adder_tree_pkg is

    type slv_vector_t is array (natural range <>) of std_logic_vector(31 downto 0); 
    
end package adder_tree_pkg;


package body adder_tree_pkg is

end package body adder_tree_pkg;